`ifndef __UART_CSR_VH__
`define __UART_CSR_VH__


`define ADDR_REG1 16'h0
`define ADDR_REG2 16'h0


`endif
