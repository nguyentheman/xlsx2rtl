`define ADDR_REG1 16'h0
`define ADDR_REG2 16'h8
